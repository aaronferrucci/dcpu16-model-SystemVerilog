typedef logic[7:0] u8;
typedef logic[15:0] u16;
typedef logic[31:0] u32;

typedef logic [3:0] t_basic_opcode;
typedef logic [5:0] t_nonbasic_opcode;
typedef logic [5:0] t_operand;

